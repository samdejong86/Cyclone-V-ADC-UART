-- lpm_pll.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity lpm_pll is
	port (
		pll_0_locked_export : out std_logic;        --  pll_0_locked.export
		pll_0_outclk0_clk   : out std_logic;        -- pll_0_outclk0.clk
		pll_0_outclk1_clk   : out std_logic;        -- pll_0_outclk1.clk
		pll_0_outclk2_clk   : out std_logic;        -- pll_0_outclk2.clk
		pll_0_outclk3_clk   : out std_logic;        -- pll_0_outclk3.clk
		pll_0_refclk_clk    : in  std_logic := '0'; --  pll_0_refclk.clk
		pll_0_reset_reset   : in  std_logic := '0'  --   pll_0_reset.reset
	);
end entity lpm_pll;

architecture rtl of lpm_pll is
	component lpm_pll_pll_0 is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			outclk_3 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component lpm_pll_pll_0;

begin

	pll_0 : component lpm_pll_pll_0
		port map (
			refclk   => pll_0_refclk_clk,    --  refclk.clk
			rst      => pll_0_reset_reset,   --   reset.reset
			outclk_0 => pll_0_outclk0_clk,   -- outclk0.clk
			outclk_1 => pll_0_outclk1_clk,   -- outclk1.clk
			outclk_2 => pll_0_outclk2_clk,   -- outclk2.clk
			outclk_3 => pll_0_outclk3_clk,   -- outclk3.clk
			locked   => pll_0_locked_export  --  locked.export
		);

end architecture rtl; -- of lpm_pll
