module controlChars(delayChar, trigSourceChar, trigSlopeChar);

output reg [7:0] delayChar  = 8'b01100100;
output reg [7:0] trigSourceChar = 8'b01110100;
output reg [7:0] trigSlopeChar = 8'b01110011;

endmodule
