module trigLevel(trigLevel);

output		    [13:0]		trigLevel = 9000;

endmodule 