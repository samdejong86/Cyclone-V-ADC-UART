module trigLevel(posTrigLevel, negTrigLevel);

output		    [13:0]		posTrigLevel = 9400;
output			 [13:0]		negTrigLevel = 7000;

endmodule 