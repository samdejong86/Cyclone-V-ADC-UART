module ExtTrigLevel(TrigSlope, TrigLevel);

output		    				TrigSlope = 1;
output			 [13:0]		TrigLevel = 10;

endmodule 