module delayVec(clk, ADC_IN, Delay);

input [13:0] ADC_IN;
input clk;


output reg [13:0] Delay [100];

always @(posedge clk) begin
   Delay[99]<=Delay[98];
   Delay[98]<=Delay[97];
   Delay[97]<=Delay[96];
   Delay[96]<=Delay[95];
   Delay[95]<=Delay[94];
   Delay[94]<=Delay[93];
   Delay[93]<=Delay[92];
   Delay[92]<=Delay[91];
   Delay[91]<=Delay[90];
   Delay[90]<=Delay[89];
   Delay[89]<=Delay[88];
   Delay[88]<=Delay[87];
   Delay[87]<=Delay[86];
   Delay[86]<=Delay[85];
   Delay[85]<=Delay[84];
   Delay[84]<=Delay[83];
   Delay[83]<=Delay[82];
   Delay[82]<=Delay[81];
   Delay[81]<=Delay[80];
   Delay[80]<=Delay[79];
   Delay[79]<=Delay[78];
   Delay[78]<=Delay[77];
   Delay[77]<=Delay[76];
   Delay[76]<=Delay[75];
   Delay[75]<=Delay[74];
   Delay[74]<=Delay[73];
   Delay[73]<=Delay[72];
   Delay[72]<=Delay[71];
   Delay[71]<=Delay[70];
   Delay[70]<=Delay[69];
   Delay[69]<=Delay[68];
   Delay[68]<=Delay[67];
   Delay[67]<=Delay[66];
   Delay[66]<=Delay[65];
   Delay[65]<=Delay[64];
   Delay[64]<=Delay[63];
   Delay[63]<=Delay[62];
   Delay[62]<=Delay[61];
   Delay[61]<=Delay[60];
   Delay[60]<=Delay[59];
   Delay[59]<=Delay[58];
   Delay[58]<=Delay[57];
   Delay[57]<=Delay[56];
   Delay[56]<=Delay[55];
   Delay[55]<=Delay[54];
   Delay[54]<=Delay[53];
   Delay[53]<=Delay[52];
   Delay[52]<=Delay[51];
   Delay[51]<=Delay[50];
   Delay[50]<=Delay[49];
   Delay[49]<=Delay[48];
   Delay[48]<=Delay[47];
   Delay[47]<=Delay[46];
   Delay[46]<=Delay[45];
   Delay[45]<=Delay[44];
   Delay[44]<=Delay[43];
   Delay[43]<=Delay[42];
   Delay[42]<=Delay[41];
   Delay[41]<=Delay[40];
   Delay[40]<=Delay[39];
   Delay[39]<=Delay[38];
   Delay[38]<=Delay[37];
   Delay[37]<=Delay[36];
   Delay[36]<=Delay[35];
   Delay[35]<=Delay[34];
   Delay[34]<=Delay[33];
   Delay[33]<=Delay[32];
   Delay[32]<=Delay[31];
   Delay[31]<=Delay[30];
   Delay[30]<=Delay[29];
   Delay[29]<=Delay[28];
   Delay[28]<=Delay[27];
   Delay[27]<=Delay[26];
   Delay[26]<=Delay[25];
   Delay[25]<=Delay[24];
   Delay[24]<=Delay[23];
   Delay[23]<=Delay[22];
   Delay[22]<=Delay[21];
   Delay[21]<=Delay[20];
   Delay[20]<=Delay[19];
   Delay[19]<=Delay[18];
   Delay[18]<=Delay[17];
   Delay[17]<=Delay[16];
   Delay[16]<=Delay[15];
   Delay[15]<=Delay[14];
   Delay[14]<=Delay[13];
   Delay[13]<=Delay[12];
   Delay[12]<=Delay[11];
   Delay[11]<=Delay[10];
   Delay[10]<=Delay[9];
   Delay[9]<=Delay[8];
   Delay[8]<=Delay[7];
   Delay[7]<=Delay[6];
   Delay[6]<=Delay[5];
   Delay[5]<=Delay[4];
   Delay[4]<=Delay[3];
   Delay[3]<=Delay[2];
   Delay[2]<=Delay[1];
   Delay[1]<=Delay[0];
	Delay[0]<=ADC_IN;
	
end

endmodule
