-- UART_pll.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity UART_pll is
	port (
		uart_pll_locked_export : out std_logic;        --  uart_pll_locked.export
		uart_pll_outclk0_clk   : out std_logic;        -- uart_pll_outclk0.clk
		uart_pll_refclk_clk    : in  std_logic := '0'; --  uart_pll_refclk.clk
		uart_pll_reset_reset   : in  std_logic := '0'  --   uart_pll_reset.reset
	);
end entity UART_pll;

architecture rtl of UART_pll is
	component UART_pll_UART_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component UART_pll_UART_pll;

begin

	uart_pll : component UART_pll_UART_pll
		port map (
			refclk   => uart_pll_refclk_clk,    --  refclk.clk
			rst      => uart_pll_reset_reset,   --   reset.reset
			outclk_0 => uart_pll_outclk0_clk,   -- outclk0.clk
			locked   => uart_pll_locked_export  --  locked.export
		);

end architecture rtl; -- of UART_pll
