
module lpm_pll (
	pll_0_locked_export,
	pll_0_outclk0_clk,
	pll_0_outclk1_clk,
	pll_0_outclk2_clk,
	pll_0_outclk3_clk,
	pll_0_refclk_clk,
	pll_0_reset_reset);	

	output		pll_0_locked_export;
	output		pll_0_outclk0_clk;
	output		pll_0_outclk1_clk;
	output		pll_0_outclk2_clk;
	output		pll_0_outclk3_clk;
	input		pll_0_refclk_clk;
	input		pll_0_reset_reset;
endmodule
