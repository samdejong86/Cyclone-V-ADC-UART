module trigLevel(trigLevel);

output		    [13:0]		trigLevel = 7000;

endmodule 